class rst_transaction extends uvm_sequence_item;
    `uvm_component_utils(rst_transaction)

    logic rst_n;

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction : new

    function string toString();
        return $sformatf("%3t - reset: %1b", $time, rst_n);
    endfunction : toString
endclass