interface reset_intf;
    logic rst;

    //get signals
    //send signals
endinterface