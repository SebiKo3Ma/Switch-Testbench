package rst_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "rst_transaction.sv"
    `include "rst_sequencer.sv"
    `include "master_driver.sv"
    `include "rst_driver.sv"
    `include "rst_monitor.sv"
    `include "rst_agent.sv"

endpackage : rst_pkg