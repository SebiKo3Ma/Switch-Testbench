package input_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "input_transaction.sv"
    `include "input_sequencer.sv"
    `include "master_driver.sv"
    `include "input_driver.sv"
    `include "input_monitor.sv"
    `include "input_agent.sv"

endpackage : input_pkg