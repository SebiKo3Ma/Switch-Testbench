package mem_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "transactions/mem_transaction.sv"
    `include "transactions/mem_write_item.sv"
    `include "transactions/mem_read_item.sv"
    `include "transactions/mem_idle_item.sv"
    `include "sequencers/mem_sequencer.sv"
    `include "drivers/mem_driver.sv"
    `include "monitors/mem_monitor.sv"
    `include "agents/mem_agent.sv"

endpackage : mem_pkg