package rst_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "transactions/rst_transaction.sv"
    `include "sequencers/rst_sequencer.sv"
    `include "drivers/rst_driver.sv"
    `include "monitors/rst_monitor.sv"
    `include "agents/rst_agent.sv"

endpackage : rst_pkg