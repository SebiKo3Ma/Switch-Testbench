interface clk_if(input clk);
endinterface