package output_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "transactions/output_transaction.sv"
    `include "sequencers/output_sequencer.sv"
    `include "drivers/output_driver.sv"
    `include "monitors/output_monitor.sv"
    `include "agents/output_agent.sv"

endpackage : output_pkg