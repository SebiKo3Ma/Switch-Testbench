package testbench_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import rst_pkg::*;
    import input_pkg::*;
    import mem_pkg::*;
    import output_pkg::*;
    `include "coverage.sv"
    `include "coverage_collector.sv"
    `include "environment.sv"
endpackage : testbench_pkg