package mem_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "mem_transaction.sv"
    `include "mem_sequencer.sv"
    `include "master_driver.sv"
    `include "mem_driver.sv"
    `include "mem_monitor.sv"
    `include "mem_agent.sv"

endpackage : mem_pkg