package testbench_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import rst_pkg::*;
    import input_pkg::*;
    import mem_pkg::*;
    import output_pkg::*;

    `include "environment.sv"
endpackage : testbench_pkg