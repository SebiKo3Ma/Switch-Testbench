package input_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "transactions/input_transaction.sv"
    `include "sequencers/input_sequencer.sv"
    `include "drivers/input_driver.sv"
    `include "monitors/input_monitor.sv"
    `include "agents/input_agent.sv"

endpackage : input_pkg