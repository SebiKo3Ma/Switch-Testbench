package input_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "input_transaction.sv"
    `include "input_if.sv"
    `include "input_sequencer.sv"
    `include "input_driver.sv"
    `include "input_monitor.sv"
    `include "input agent.sv"

endpackage : input_pkg