package rst_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "rst_transaction.sv"
    `include "clk_rst_if.sv"
    `include "rst_sequencer.sv"
    `include "rst_driver.sv"
    `include "rst_monitor.sv"
    `include "rst agent.sv"

endpackage : rst_pkg