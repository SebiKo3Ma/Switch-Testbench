interface clk_intf(input clk);
    logic clk;
    
    //get signals
    //send signals
endinterface