interface output_intf;
    logic [7:0] port_out;   //serial 1-byte data output
    logic       port_ready; //ready signal for data output
    logic       port_read;  //read input signal for output port

    //get signals
    //send signals
endinterface